`define SUPPORT_RV32C 1
`define SUPPORT_RV32M 1
`define ENABLE_COUNTERS 1
`define ENABLE_IRQ 1
`define ENABLE_TIMER 1
`define TWO_STAGE_SHIFT 1
`define TWO_CYCLE_COMPARE 0
`define TWO_CYCLE_ALU 0
`define BARREL_SHIFTER 0
`define CATCH_MISALIGN 1
`define CATCH_ILLINSN 1
`define ENABLE_DEBUG
`define I_MEM_K_BYTE 8
`define BUILD_LOAD
`define SW_BIN_PATH "F:/code/fpga/MIC_HDMI_FINISHED/ram32.hex"
`define D_MEM_K_BYTE 8
`define ENABLE_HSP 0
`define HSP_VALUE_DEF 32'h0
`define ENABLE_OPEN_AHB
`define ENABLE_WB_UART
